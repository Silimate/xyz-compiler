module _ONE_(Y);
	output wire Y = 1;
endmodule
module _ZERO_(Y);
	output wire Y = 0;
endmodule
